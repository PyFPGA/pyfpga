`define DEFAULT_FREQ 25000000
`define DEFAULT_SECS 1
