`define INCLUDE
