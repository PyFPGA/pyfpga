entity Top1 is
end entity Top1;

-- entity Top2 is
-- end entity Top1;
