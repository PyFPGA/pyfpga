`define INCLUDE2
