`define DEFAULT_FREQ 25000000
