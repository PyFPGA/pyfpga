`define DEFAULT_SECS 1
