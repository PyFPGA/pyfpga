`define INCLUDE1
