../../hdl/blinking.vhdl